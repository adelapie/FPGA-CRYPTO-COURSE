
-- Copyright (c) 2013 Antonio de la Piedra

-- This program is free software: you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.

-- This program is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.

-- You should have received a copy of the GNU General Public License
-- along with this program.  If not, see <http://www.gnu.org/licenses/>.

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
  
ENTITY tb_round_f IS
END tb_round_f;
 
ARCHITECTURE behavior OF tb_round_f IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT round_f
    PORT(clk : in std_logic;
	      rst : in std_logic;
         enc : in std_logic;
         rc_in : IN  std_logic_vector(31 downto 0);
         a_0_in : IN  std_logic_vector(31 downto 0);
         a_1_in : IN  std_logic_vector(31 downto 0);
         a_2_in : IN  std_logic_vector(31 downto 0);
         a_3_in : IN  std_logic_vector(31 downto 0);
         k_0_in : IN  std_logic_vector(31 downto 0);
         k_1_in : IN  std_logic_vector(31 downto 0);
         k_2_in : IN  std_logic_vector(31 downto 0);
         k_3_in : IN  std_logic_vector(31 downto 0);
         a_0_out : OUT  std_logic_vector(31 downto 0);
         a_1_out : OUT  std_logic_vector(31 downto 0);
         a_2_out : OUT  std_logic_vector(31 downto 0);
         a_3_out : OUT  std_logic_vector(31 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
	signal enc : std_logic := '0';
	signal rst : std_logic := '0';

   signal rc_in : std_logic_vector(31 downto 0) := (others => '0');
   signal a_0_in : std_logic_vector(31 downto 0) := (others => '0');
   signal a_1_in : std_logic_vector(31 downto 0) := (others => '0');
   signal a_2_in : std_logic_vector(31 downto 0) := (others => '0');
   signal a_3_in : std_logic_vector(31 downto 0) := (others => '0');
   signal k_0_in : std_logic_vector(31 downto 0) := (others => '0');
   signal k_1_in : std_logic_vector(31 downto 0) := (others => '0');
   signal k_2_in : std_logic_vector(31 downto 0) := (others => '0');
   signal k_3_in : std_logic_vector(31 downto 0) := (others => '0');

 	--Outputs
   signal a_0_out : std_logic_vector(31 downto 0);
   signal a_1_out : std_logic_vector(31 downto 0);
   signal a_2_out : std_logic_vector(31 downto 0);
   signal a_3_out : std_logic_vector(31 downto 0);

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: round_f PORT MAP (
			 clk => clk,
			 rst => rst,
          enc => enc,
          rc_in => rc_in,
          a_0_in => a_0_in,
          a_1_in => a_1_in,
          a_2_in => a_2_in,
          a_3_in => a_3_in,
          k_0_in => k_0_in,
          k_1_in => k_1_in,
          k_2_in => k_2_in,
          k_3_in => k_3_in,
          a_0_out => a_0_out,
          a_1_out => a_1_out,
          a_2_out => a_2_out,
          a_3_out => a_3_out
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
		wait for clk_period + clk_period/2;
		rst <= '1';
		wait for clk_period;
		rst <= '0';
		
		rc_in  <= X"00000080";
		
		a_0_in <= X"61396c93";
		a_1_in <= X"637434b8";		
		a_2_in <= X"fc6559a9";
		a_3_in <= X"5b643f2c";

		k_0_in <= X"1c1c1c1c";
		k_1_in <= X"1c1c1c1c";
		k_2_in <= X"1c1c1c1c";
		k_3_in <= X"1c1c1c1c";

		wait for clk_period;

--		assert a_0_out = X"febb00d0"
--			report "ROUND ERROR (a_0)" severity FAILURE;		
--			
--		assert a_1_out = X"074ee42e"
--			report "ROUND ERROR (a_1)" severity FAILURE;		
--
--		assert a_2_out = X"dde647ab"
--			report "ROUND ERROR (a_2)" severity FAILURE;		
--			
--		assert a_3_out = X"3207ef78"
--			report "ROUND ERROR (a_3)" severity FAILURE;			
			
      wait;
   end process;

END;
